class i2cmb_random_transaction_test extends i2cmb_test_base;


  function new(string name = "", ncsu_component_base parent = null); 
    super.new(name,parent);
    
  endfunction

endclass
